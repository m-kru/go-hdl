--thdl:ignore
clk_20_i => clk_40_i

   --thdl:ignore
   clk_50 => clk_70
