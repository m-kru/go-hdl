clk_20_i => clk_40_i --hdl:ignore  

   if rst_p = '0' then --hdl:ignore
