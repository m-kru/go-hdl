--hdl:ignore
clk_20_i => clk_40_i

   --hdl:ignore
   clk_50 => clk_70
