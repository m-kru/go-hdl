clk_20_i => clk_40_i --thdl:ignore  

   if rst_p = '0' then --thdl:ignore
