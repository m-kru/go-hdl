process (clk_i)
begin
  if (rising_edge(clk_i)) then
  end if;
end process;
