process (foo) is
   if rising_edge(bar) then
   end if;
begin
end process;
