process (tx_clk(1))
begin
  if rising_edge(tx_clk(1)) then
    end if;
  end if;
end process;
