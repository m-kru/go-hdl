process is
   if rising_edge(clk) then
   end if;
begin
end process;
